module Top(
    // q90weqw09didlausd
);
endmodule